library verilog;
use verilog.vl_types.all;
entity Fred_testbench is
end Fred_testbench;
