library verilog;
use verilog.vl_types.all;
entity nordstrom_testbench is
end nordstrom_testbench;
