library verilog;
use verilog.vl_types.all;
entity last2Digits_testbench is
end last2Digits_testbench;
